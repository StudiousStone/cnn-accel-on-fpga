/*
* Created           : cheng liu
* Date              : 2016-04-26
*
* Description:
* 
* Verify the read master port and write master port 
* 
* 
*/

`timescale 1ns/1ns

module avlon_tb;

parameter CLK_PERIOD = 10;
parameter DATA_SIZE = 1024;
parameter TILE_SIZE = 128;
parameter R_PORT = 1;
parameter W_PORT = 1;

localparam AW = 12;
localparam DW = 32;
localparam CW = 8;
localparam RES = 24;
localparam XAW = 32;
localparam XDW = 128;
localparam WCNT =(XDW/DW);

wire  [R_PORT-1:0]        rmst_fixed_location;   // fixed_location
wire  [R_PORT*XAW-1:0]    rmst_read_base;        // read_base
wire  [R_PORT*XAW-1:0]    rmst_read_length;      // read_length
wire  [R_PORT*CW-1: 0]    rmst_read_length_tmp;
wire  [R_PORT-1:0]        rmst_go;               // go
wire  [R_PORT-1:0]        rmst_done;             // done
wire  [R_PORT-1:0]        rmst_user_read_buffer;      // read_buffer
wire  [R_PORT*128-1:0]    rmst_user_buffer_data;      // buffer_output_data
wire  [R_PORT-1:0]        rmst_user_data_available;   // data_available

wire  [W_PORT-1:0]        wmst_fixed_location;   // fixed_location
wire  [W_PORT*XAW-1:0]    wmst_write_base;       // write_base
wire  [W_PORT*XAW-1:0]    wmst_write_length;     // write_length
wire  [W_PORT*CW-1: 0]    wmst_write_length_tmp;
wire  [W_PORT-1:0]        wmst_go;               // go
wire  [W_PORT-1:0]        wmst_done;             // done
wire  [W_PORT-1:0]        wmst_user_write_buffer;// write_buffer
wire  [W_PORT*128-1:0]    wmst_user_write_data;  // buffer_input_data
wire  [W_PORT-1:0]        wmst_user_buffer_full;      

reg                       config_start;
wire                      config_done;

wire            [DW-1: 0] param_raddr;
wire            [DW-1: 0] param_waddr;
wire            [AW-1: 0] param_iolen;

wire                      load_data_start;
wire                      load_data_done;
wire                      store_data_start;
wire                      store_data_done;

//wire                      rmst_wr_ena;
//wire            [DW-1: 0] rmst_wr_data;
//wire            [AW-1: 0] rmst_wr_addr;

//wire            [AW-1: 0] wmst_rd_addr;
//wire            [DW-1: 0] wmst_rd_data;

wire            [DW-1: 0] rmst_load_data;
wire                      load_fifo_push;
wire                      load_fifo_almost_full;

wire            [DW-1: 0] wmst_store_data;
wire                      store_fifo_pop;
wire                      store_fifo_empty;

reg         clk = 0;
reg         rst = 0;
wire        task_done;

always # (CLK_PERIOD / 2) clk = ~clk;

initial begin
    rst = 1;
    config_start <= 1'b0;

    repeat (5) begin
        @(posedge clk);
    end
    rst = 0; 

    @(posedge clk)
    config_start <= 1'b1;

    @(posedge clk)
    config_start <= 1'b0;

end

transfer_config #(
    .AW (AW),  // Internal memory address width
    .DW (DW),  // Internal data width
    .CW (CW),  // maxium number of configuration paramters is (2^CW).
    .DATA_SIZE (DATA_SIZE)
)transfer_config(
    .config_start (config_start),
    .config_done  (config_done), 

    .param_raddr  (param_raddr),
    .param_waddr  (param_waddr),
    .param_iolen  (param_iolen),

    .task_done    (task_done), // computing task is done. (original name: flag_over)
    .store_data_done (store_data_done),
    
    .rst          (rst),
    .clk          (clk)
);


sig_delay #(
    .D (10)
) sig_delay0 (
    .sig_in (config_done),
    .sig_out (load_data_start),

    .clk (clk),
    .rst (rst)
);


sig_delay #(
    .D (10)
) sig_delay (
    .sig_in (load_data_start),
    .sig_out (store_data_start),

    .clk (clk),
    .rst (rst)
);

rmst_to_fifo_tile #(
    .AW (AW),
    .CW (CW),
    .DW (DW),
    .XAW (XAW),
    .XDW (XDW)
) rmst_in_fm (
    .param_raddr           (param_raddr),
    .param_iolen           (param_iolen),
    .config_done           (config_done),

    .rmst_fixed_location   (rmst_fixed_location),
    .rmst_read_base        (rmst_read_base),
    .rmst_read_length      (rmst_read_length_tmp),
    .rmst_go               (rmst_go),
    .rmst_done             (rmst_done),

    .rmst_user_read_buffer (rmst_user_read_buffer),
    .rmst_user_buffer_data (rmst_user_buffer_data),
    .rmst_user_data_available (rmst_user_data_available),

    //.rmst_wr_ena              (rmst_wr_ena),
    //.rmst_wr_data             (rmst_wr_data),
    //.rmst_wr_addr             (rmst_wr_addr),

    .load_data_done           (load_data_done),
    .load_data_start          (load_data_start),

    .rmst_load_data           (rmst_load_data),
    .load_fifo_push           (load_fifo_push),
    .load_fifo_almost_full    (load_fifo_almost_full),

    .clk                   (clk),
    .rst                   (rst)
);

wmst_to_fifo_tile #(
    .AW (AW),
    .CW (CW),
    .DW (DW),
    .XAW (XAW),
    .XDW (XDW)
) wmst_out_fm (
    .param_waddr           (param_waddr),
    .param_iolen           (param_iolen),
    .config_done           (config_done),
    
    .wmst_fixed_location   (wmst_fixed_location),
    .wmst_write_base       (wmst_write_base),
    .wmst_write_length     (wmst_write_length_tmp),
    .wmst_go               (wmst_go),
    .wmst_done             (wmst_done),

    .wmst_user_write_buffer(wmst_user_write_buffer),
    .wmst_user_write_data  (wmst_user_write_data),
    .wmst_user_buffer_full (wmst_user_buffer_full),

    .store_data_done       (store_data_done),
    .store_data_start      (store_data_start),

    //.wmst_rd_data          (wmst_rd_data),
    //.wmst_rd_addr          (wmst_rd_addr),

    .wmst_store_data       (wmst_store_data),
    .store_fifo_pop        (store_fifo_pop),
    .store_fifo_empty      (store_fifo_empty),
    
    .clk                   (clk),
    .rst                   (rst)
);

assign rmst_read_length = {24'b0, rmst_read_length_tmp};
assign wmst_write_length = {24'b0, wmst_write_length_tmp};

mem_top #(
    .R_PORT (R_PORT),
    .W_PORT (W_PORT)
) mem_model(
    .read_control_fixed_location  (rmst_fixed_location),
    .read_control_read_base       (rmst_read_base),
    .read_control_read_length     (rmst_read_length),
    .read_control_go              (rmst_go), 
    .read_control_done            (rmst_done), 
    .read_user_read_buffer        (rmst_user_read_buffer),
    .read_user_buffer_output_data (rmst_user_buffer_data),
    .read_user_data_available     (rmst_user_data_available),

    .write_control_fixed_location (wmst_fixed_location),
    .write_control_write_base     (wmst_write_base),
    .write_control_write_length   (wmst_write_length),
    .write_control_go             (wmst_go),
    .write_control_done           (wmst_done), 
    .write_user_write_buffer      (wmst_user_write_buffer),
    .write_user_buffer_input_data (wmst_user_write_data),
    .write_user_buffer_full       (wmst_user_buffer_full), 
    
    .clk (clk),
    .rst (rst)
);

/*
 dp_mem #(      .AW(AW),      .DW(DW),      .DATA_SIZE (DATA_SIZE)
  ) dp_mem (
      .clk (clk),
      .rst (rst),
      .data_in (rmst_wr_data),
      .raddr (wmst_rd_addr),
      .waddr (rmst_wr_addr),
      .wena (rmst_wr_ena),
      .data_out (wmst_rd_data)
  );
*/


scfifo	SCFF (
    .aclr           (rst),
    .clock          (clk),
    .data           (rmst_load_data),
    .rdreq          (store_fifo_pop),
    .sclr           (1'b0),
    .wrreq          (load_fifo_push),
    .almost_empty   (),
    .almost_full    (load_fifo_almost_full),
    .empty          (store_fifo_empty),
    .full           (),
    .q              (wmst_store_data),
    .usedw          (),
    .eccstatus ());
defparam
    SCFF.add_ram_output_register = "OFF",
    SCFF.almost_empty_value = 8,
    SCFF.almost_full_value = 250,
    SCFF.intended_device_family = "Cyclone V",
    SCFF.lpm_hint = "RAM_BLOCK_TYPE=M10K",
    SCFF.lpm_numwords = 256,
    SCFF.lpm_showahead = "OFF",
    SCFF.lpm_type = "scfifo",
    SCFF.lpm_width = 32,
    SCFF.lpm_widthu = 8,
    SCFF.overflow_checking = "ON",
    SCFF.underflow_checking = "ON",
    SCFF.use_eab = "ON";


endmodule
