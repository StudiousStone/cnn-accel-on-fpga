/*
* Created           : cheng liu
* Date              : 2016-04-26
*
* Description:
* 
* Verify the read master port and write master port 
* 
* 
*/

`timescale 1ns/1ns

module avlon_tb;

parameter CLK_PERIOD = 10;
parameter R_PORT = 1;
parameter W_PORT = 1;

parameter AW = 12;
parameter CW = 16;
parameter DW = 32;
parameter XAW = 32;
parameter XDW = 128;
    parameter N = 16;
    parameter M = 16;
    parameter R = 32;
    parameter C = 16;
    parameter Tn = 8;
    parameter Tm = 8;
    parameter Tr = 16;
    parameter Tc = 8;
parameter S = 1;
parameter K = 3;

localparam WCNT =(XDW/DW);

wire  [R_PORT-1:0]        rmst_fixed_location;   // fixed_location
wire  [R_PORT*XAW-1:0]    rmst_read_base;        // read_base
wire  [R_PORT*XAW-1:0]    rmst_read_length;      // read_length
wire  [R_PORT*CW-1: 0]    rmst_read_length_tmp;
wire  [R_PORT-1:0]        rmst_go;               // go
wire  [R_PORT-1:0]        rmst_done;             // done
wire  [R_PORT-1:0]        rmst_user_read_buffer;      // read_buffer
wire  [R_PORT*128-1:0]    rmst_user_buffer_data;      // buffer_output_data
wire  [R_PORT-1:0]        rmst_user_data_available;   // data_available

wire  [W_PORT-1:0]        wmst_fixed_location;   // fixed_location
wire  [W_PORT*XAW-1:0]    wmst_write_base;       // write_base
wire  [W_PORT*XAW-1:0]    wmst_write_length;     // write_length
wire  [W_PORT*CW-1: 0]    wmst_write_length_tmp;
wire  [W_PORT-1:0]        wmst_go;               // go
wire  [W_PORT-1:0]        wmst_done;             // done
wire  [W_PORT-1:0]        wmst_user_write_buffer;// write_buffer
wire  [W_PORT*128-1:0]    wmst_user_write_data;  // buffer_input_data
wire  [W_PORT-1:0]        wmst_user_buffer_full;      

reg                       load_start;
wire                      load_done;
reg                       store_start;
wire                      store_done;

wire            [DW-1: 0] rmst_load_data;
wire                      load_fifo_push;
wire                      load_fifo_almost_full;

wire            [DW-1: 0] wmst_store_data;
wire                      store_fifo_pop;
wire                      store_fifo_empty;

reg             [CW-1: 0] tile_base_m;
reg             [CW-1: 0] tile_base_row;
reg             [CW-1: 0] tile_base_col;

reg         clk = 0;
reg         rst = 0;

always # (CLK_PERIOD / 2) clk = ~clk;

initial begin
    rst = 1;
    load_start <= 1'b0;
    store_start <= 1'b0;

    tile_base_m = 0;
    tile_base_row = 0;
    tile_base_col = 0;

    repeat (5) begin
        @(posedge clk);
    end
    rst = 0; 

    @(posedge clk)
    load_start <= 1'b1;

    @(posedge clk)
    load_start <= 1'b0;

    repeat (10) begin
        @(posedge clk);
    end
    store_start <= 1'b1;

    @(posedge clk)
    store_start <= 1'b0;

end

rmst_to_fifo_tile #(
    .AW (AW),
    .CW (CW),
    .DW (DW),
    .XAW (XAW),
    .XDW (XDW),
        .N (N),
        .M (M),
        .R (R),
        .C (C),
        .Tn (Tn),
        .Tm (Tm),
        .Tr (Tr),
        .Tc (Tc),
        .S (S),
        .K (K)
) rmst_in_fm (
    .rmst_fixed_location   (rmst_fixed_location),
    .rmst_read_base        (rmst_read_base),
    .rmst_read_length      (rmst_read_length_tmp),
    .rmst_go               (rmst_go),
    .rmst_done             (rmst_done),

    .rmst_user_read_buffer (rmst_user_read_buffer),
    .rmst_user_buffer_data (rmst_user_buffer_data),
    .rmst_user_data_available (rmst_user_data_available),

    .load_done             (load_done),
    .load_start            (load_start),

    .rmst_load_data           (rmst_load_data),
    .load_fifo_push           (load_fifo_push),
    .load_fifo_almost_full    (load_fifo_almost_full),

    .tile_base_m (tile_base_m),
    .tile_base_row (tile_base_row),
    .tile_base_col (tile_base_col),

    .clk                   (clk),
    .rst                   (rst)
);

wmst_to_fifo_tile #(
    .AW (AW),
    .CW (CW),
    .DW (DW),
    .XAW (XAW),
    .XDW (XDW),
        .N (N),
        .M (M),
        .R (R),
        .C (C),
        .Tn (Tn),
        .Tm (Tm),
        .Tr (Tr),
        .Tc (Tc),
        .S (S),
        .K (K)
) wmst_out_fm (
    .wmst_fixed_location   (wmst_fixed_location),
    .wmst_write_base       (wmst_write_base),
    .wmst_write_length     (wmst_write_length_tmp),
    .wmst_go               (wmst_go),
    .wmst_done             (wmst_done),

    .wmst_user_write_buffer(wmst_user_write_buffer),
    .wmst_user_write_data  (wmst_user_write_data),
    .wmst_user_buffer_full (wmst_user_buffer_full),

    .store_done       (store_done),
    .store_start      (store_start),

    .wmst_store_data       (wmst_store_data),
    .store_fifo_pop        (store_fifo_pop),
    .store_fifo_empty      (store_fifo_empty),

    .tile_base_m (tile_base_m),
    .tile_base_row (tile_base_row),
    .tile_base_col (tile_base_col),
    
    .clk                   (clk),
    .rst                   (rst)
);

assign rmst_read_length = {16'b0, rmst_read_length_tmp};
assign wmst_write_length = {16'b0, wmst_write_length_tmp};

mem_top #(
    .R_PORT (R_PORT),
    .W_PORT (W_PORT)
) mem_model(
    .read_control_fixed_location  (rmst_fixed_location),
    .read_control_read_base       (rmst_read_base),
    .read_control_read_length     (rmst_read_length),
    .read_control_go              (rmst_go), 
    .read_control_done            (rmst_done), 
    .read_user_read_buffer        (rmst_user_read_buffer),
    .read_user_buffer_output_data (rmst_user_buffer_data),
    .read_user_data_available     (rmst_user_data_available),

    .write_control_fixed_location (wmst_fixed_location),
    .write_control_write_base     (wmst_write_base),
    .write_control_write_length   (wmst_write_length),
    .write_control_go             (wmst_go),
    .write_control_done           (wmst_done), 
    .write_user_write_buffer      (wmst_user_write_buffer),
    .write_user_buffer_input_data (wmst_user_write_data),
    .write_user_buffer_full       (wmst_user_buffer_full), 
    
    .clk (clk),
    .rst (rst)
);

scfifo	SCFF (
    .aclr           (rst),
    .clock          (clk),
    .data           (rmst_load_data),
    .rdreq          (store_fifo_pop),
    .sclr           (1'b0),
    .wrreq          (load_fifo_push),
    .almost_empty   (),
    .almost_full    (load_fifo_almost_full),
    .empty          (store_fifo_empty),
    .full           (),
    .q              (wmst_store_data),
    .usedw          (),
    .eccstatus ());
defparam
    SCFF.add_ram_output_register = "OFF",
    SCFF.almost_empty_value = 8,
    SCFF.almost_full_value = 250,
    SCFF.intended_device_family = "Cyclone V",
    SCFF.lpm_hint = "RAM_BLOCK_TYPE=M10K",
    SCFF.lpm_numwords = 256,
    SCFF.lpm_showahead = "OFF",
    SCFF.lpm_type = "scfifo",
    SCFF.lpm_width = 32,
    SCFF.lpm_widthu = 8,
    SCFF.overflow_checking = "ON",
    SCFF.underflow_checking = "ON",
    SCFF.use_eab = "ON";


endmodule
