/*
* Created           : Cheng Liu 
* Date              : 2016-04-25
*
* Description:
* This is a simple dual port memory allowing both read and write 
* operations at the same time as long as there are no read/write 
* conflicts. Note that the read port and write port are shared between 
* the internal softmax computing logic and the external system bus.

softmax_dp_mem #(
    .AW (),
    .DW (),
    .XAW (),
    .XDW (),
    .WCNT ()

)(
    // Port connected to the read master
    .rmst_fixed_location (),
    .rmst_read_base (),
    .rmst_read_length (),
    .rmst_go (),
    .rmst_done (),

    .rmst_user_read_buffer (),
    .rmst_user_buffer_data (),
    .rmst_user_data_available (), 

    // Port connected to the write master
    .wmst_fixed_location (),
    .wmst_write_base (),
    .wmst_write_length (),
    .wmst_go (),
    .wmst_done (),
    .wmst_user_write_data (),
    .wmst_user_write_buffer (),
    .wmst_user_buffer_full (),

    // Parameters from the configuration module
    .param_raddr (),
    .param_iolen (),
    .param_waddr (),

    .load_data_done (),
    .store_data_done (),

    // Internal memomry port to the softmax_core
    .internal_wr_addr (),
    .internal_wr_data (),
    .internal_wr_ena (),

    .internal_rd_addr (),
    .internal_rd_data (),

    .store_data_start (),
    .load_data_start (),

    .rst (),
    .clk ()
);

*/

// synposys translate_off
`timescale 1ns/100ps
// synposys translate_on

module softmax_dp_mem #(
    parameter AW = 12,
    parameter DW = 32,
    parameter XAW = 32,
    parameter XDW = 128

)(
    // Port connected to the read master
    output                             rmst_fixed_location,
    output                   [XAW-1:0] rmst_read_base,
    output                   [XAW-1:0] rmst_read_length,
    output                             rmst_go,
    input                              rmst_done,

    output                             rmst_user_read_buffer,
    input                    [XDW-1:0] rmst_user_buffer_data,
    input                              rmst_user_data_available, 

    // Port connected to the write master
    output                             wmst_fixed_location,
    output                  [XAW-1: 0] wmst_write_base,
    output                  [XAW-1: 0] wmst_write_length,
    output                             wmst_go,
    input                              wmst_done,
    output                  [XDW-1: 0] wmst_user_write_data,
    output                             wmst_user_write_buffer,
    input                              wmst_user_buffer_full,

    // Parameters from the configuration module
    input                   [XAW-1: 0] param_raddr,
    input                    [AW-1: 0] param_iolen,
    input                   [XAW-1: 0] param_waddr,

    output                             load_data_done,
    output                             store_data_done,

    // Internal memomry port to the softmax_core
    input                    [AW-1: 0] internal_wr_addr,
    input                    [DW-1: 0] internal_wr_data,
    input                              internal_wr_ena,

    input                    [AW-1: 0] internal_rd_addr,
    output                   [DW-1: 0] internal_rd_data,

    input                              store_data_start,
    input                              load_data_start,

    input                              rst,
    input                              clk
);

    localparam WCNT = (XDW/DW);
    // Internal memory port to the read master
    wire                     [AW-1: 0] rmst_wr_addr;
    wire                     [DW-1: 0] rmst_wr_data;
    wire                               rmst_wr_ena;

    // Internal memory port to the write master
    wire                     [AW-1: 0] wmst_rd_addr;
    wire                     [DW-1: 0] wmst_rd_data;
    wire                               load_data_start_d1;

    reg                     [XAW-1: 0] raddr;
    reg                     [XAW-1: 0] waddr;
    reg                      [AW-1: 0] iolen;
    reg                      [AW-1: 0] rmst_cnt;
    reg                      [AW-1: 0] wmst_cnt;
    reg                     [XDW-1: 0] rmst_rd_data;
    reg                    [WCNT-1: 0] rmst_word_ena;
    reg                    [WCNT-1: 0] wmst_word_ena;

    reg                     [XDW-1: 0] write_buffer_data_reg;
    wire                   [WCNT-1: 0] rmst_word_ena_d1;
    wire                   [WCNT-1: 0] wmst_word_ena_d2;
    wire                   [WCNT-1: 0] rmst_word_ena_d2;

    // Lock the parameters
    always@(posedge clk) begin
        if(rst == 1'b1) begin
            raddr <= 0;
            waddr <= 0;
            iolen <= 0;
        end
        else if(load_data_start == 1'b1) begin
            raddr <= param_raddr;
            waddr <= param_waddr;
            iolen <= param_iolen;
        end
        else begin
            raddr <= raddr;
            waddr <= waddr;
            iolen <= iolen; 
        end
    end

    sig_delay #(
        .D (WCNT)
    ) sig_delay1 (
        .sig_in (rmst_done),
        .sig_out (load_data_done),

        .clk (clk),
        .rst (rst)
    );

    assign rmst_fixed_location = 1'b0;
    assign rmst_read_base = raddr;
    assign rmst_read_length = iolen << 2;

    always@(posedge clk or posedge rst) begin
        if(rst == 1'b1) begin
            rmst_word_ena <= 0;
        end
        else if(rmst_user_data_available == 1'b1 && (rmst_word_ena[WCNT-1] == 1'b1 || rmst_word_ena == 0)) begin
            rmst_word_ena <= 1;
        end
        else if(rmst_user_data_available == 1'b0 && rmst_word_ena[WCNT-1] == 1'b1) begin
            rmst_word_ena <= 0;
        end
        else begin
            rmst_word_ena <= {rmst_word_ena[WCNT-2: 0], rmst_word_ena[WCNT-1]};
        end
    end

    data_delay #(
        .D (1),
        .DW (WCNT)
    ) data_delay0 (
        .clk (clk),        
        .data_in (rmst_word_ena),
        .data_out (rmst_word_ena_d1)
    );
    
    data_delay #(
        .D (1),
        .DW (WCNT)
    ) data_delay1 (
        .clk (clk),        
        .data_in (rmst_word_ena_d1),
        .data_out (rmst_word_ena_d2)
    );

    // The test bench may be wrong. The read buffer signal behaves as a read request.
    // It guess it may take XDW as the data pop granularity from the Avlon interface FIFO.
    assign rmst_user_read_buffer = rmst_user_data_available && (|rmst_word_ena)[WCNT-1]; 
    //assign rmst_user_read_buffer = rmst_user_data_available && (|rmst_word_ena); 
    always@(posedge clk or posedge rst) begin
        if(rst == 1'b1) begin
            rmst_rd_data <= 0;
        end
        else if(rmst_user_data_available == 1'b1 && rmst_word_ena_d1[0] == 1'b1) begin
            rmst_rd_data <= rmst_user_buffer_data;
        end
        else begin
            rmst_rd_data <= {32'b0, rmst_rd_data[XDW-1: 32]};
        end
    end

    assign rmst_wr_data = rmst_rd_data[31: 0];
    assign rmst_wr_ena = |rmst_word_ena_d2;
    assign rmst_wr_addr = rmst_cnt;

    // Generate rd address for internal memory write port.
    always@(posedge clk or posedge rst) begin
        if(rst == 1'b1) begin
            rmst_cnt <= 0;
        end
        else if(rmst_wr_ena == 1'b1) begin
            rmst_cnt <= rmst_cnt + 1;
        end
        else begin // clear memory for future writing iteration
            rmst_cnt <= 0;
        end
    end

    assign wmst_fixed_location = 1'b0;
    assign wmst_write_base = waddr;
    assign wmst_write_length = iolen << 2; 

    always@(posedge clk or posedge rst) begin
        if(rst == 1'b1) begin
            wmst_word_ena <= 0;
        end
        else if(store_data_start == 1'b1 && wmst_user_buffer_full == 1'b0) begin
            wmst_word_ena <= 1;
        end
        else if(wmst_user_buffer_full == 1'b1) begin
            wmst_word_ena <= wmst_word_ena;
        end
        else if(wmst_cnt == (iolen-1)) begin
            wmst_word_ena <= 0;
        end
        else begin
            wmst_word_ena <= {wmst_word_ena[WCNT-2: 0], wmst_word_ena[WCNT-1]};
        end
    end

    reg                                write_buffer_reg;
    always@(posedge clk or posedge rst) begin
        if(rst == 1'b1) begin
            write_buffer_reg <= 1'b0;
        end
        else if(wmst_word_ena_d2[WCNT-1] == 1'b1 && wmst_user_buffer_full == 1'b0) begin
            write_buffer_reg <= 1'b1;
        end
        else begin
            write_buffer_reg <= 1'b0;
        end
    end
    
    assign wmst_user_write_buffer = write_buffer_reg;

    always@(posedge clk or posedge rst) begin
        if(rst == 1'b1) begin
            wmst_cnt <= 0;
        end
        else if(store_data_start == 1'b1 && wmst_user_buffer_full == 1'b0) begin
            wmst_cnt <= 0;
        end
        else if(((|wmst_word_ena) == 1'b1) && wmst_user_buffer_full == 1'b0) begin
            wmst_cnt <= wmst_cnt + 1;
        end
        else if((wmst_word_ena[WCNT-1] == 1'b1 && wmst_user_buffer_full == 1'b1)) begin
            wmst_cnt <= wmst_cnt;
        end
        else if(wmst_cnt == (iolen-1)) begin
            wmst_cnt <= 0;
        end
        else begin
            wmst_cnt <= wmst_cnt;
        end
    end

    // Write transmission starts when the first 128bit data is ready
    reg                                go_reg;
    always@(posedge clk or posedge rst) begin
        if(rst == 1'b1) begin
            go_reg <= 1'b0;
        end
        else if(wmst_cnt == 4) begin
            go_reg <= 1'b1;
        end
        else begin
            go_reg <= 1'b0;
        end
    end
    
    sig_delay #(
        .D (1)
    ) sig_delay2 (
        .sig_in (go_reg),
        .sig_out (wmst_go),

        .clk (clk),
        .rst (rst)
    );
    
    data_delay #(
        .D (2),
        .DW (WCNT)
    ) data_delay2 (
        .clk (clk),        
        .data_in (wmst_word_ena),
        .data_out (wmst_word_ena_d2)
    );
   
    always@(posedge clk or posedge rst) begin
        if(rst == 1'b1) begin
            write_buffer_data_reg <= 0;
        end
        else if((|wmst_word_ena_d2) == 1'b1) begin
            write_buffer_data_reg <= {wmst_rd_data, write_buffer_data_reg[XDW-1: 32]};
        end
        else begin
            write_buffer_data_reg <= write_buffer_data_reg;
        end
    end

    assign wmst_user_write_data = write_buffer_data_reg;

    assign wmst_rd_addr = wmst_cnt;

    // Assume that write operation starts WAR_DELAY cycles later
    sig_delay #(
        .D (1)
    ) sig_delay3 (
        .sig_in (load_data_start,
        .sig_out (load_data_start_d1),

        .clk (clk),
        .rst (rst)
    );
    
    /*
    sig_delay #(
        .D (RAW_DELAY)
    ) sig_delay4 (
        .sig_in (config_done),
        .sig_out (load_data_start),

        .clk (clk),
        .rst (rst)
    );
    */

    assign rmst_go = load_data_start_d1;

    assign store_data_done = wmst_done;

    wire                               wr_ena;
    wire                     [AW-1: 0] wr_addr;
    wire                     [DW-1: 0] wr_data;
    wire                     [AW-1: 0] rd_addr;
    wire                     [DW-1: 0] rd_data;
    reg                                wr_sel;
    reg                                rd_sel;

    always@(posedge clk or posedge rst) begin
        if(rst == 1'b1) begin
            wr_sel <= 1'b0;
        end
        else if(load_data_start == 1'b1) begin
            wr_sel <= 1'b1;
        end
        else if(load_data_done == 1'b1) begin
            wr_sel <= 1'b0;
        end
    end

    always@(posedge clk or posedge rst) begin
        if(rst == 1'b1) begin
            rd_sel <= 1'b0;
        end
        else if(store_data_start == 1'b1) begin
            rd_sel <= 1'b1;
        end
        else if(store_data_done == 1'b1) begin
            rd_sel <= 1'b0;
        end
    end

    assign wr_data = wr_sel ? rmst_wr_data : internal_wr_data;
    assign wr_ena = wr_sel ? rmst_wr_ena : internal_wr_ena;
    assign wr_addr = wr_sel ? rmst_wr_addr : internal_wr_addr;
    assign rd_addr = rd_sel ? wmst_rd_addr : internal_rd_addr;
    assign wmst_rd_data = rd_sel ? rd_data : 0;
    assign internal_rd_data = rd_sel ? 0 : rd_data;
    
    dp_mem #(
        .AW(AW),
        .DW(DW)
    ) dp_mem (
        .clk (clk),
        .rst (rst),
        .data_in (wr_data),
        .raddr (rd_addr),
        .waddr (wr_addr),
        .wena (wr_ena),
        .data_out (rd_data)
    );

endmodule

